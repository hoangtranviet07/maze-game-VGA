--Package statements
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
entity sevseg is 
port(SW  : in STD_LOGIC_VECTOR(7 downto 0);
	  HEX0, HEX1: out STD_LOGIC_VECTOR(0 to 6));
end entity; 
architecture decoder_arch of sevseg is 
	begin 
	with (SW) select 
	 HEX0 <= "0000001" when "00000000", -- 0 
					"1001111" when "00000001", -- 1
					"0010010" when "00000010", -- 2
					"0000110" when "00000011", -- 3
					"1001100" when "00000100", -- 4
					"0100100" when "00000101", -- 5
					"0100000" when "00000110", -- 6 
					"0001111" when "00000111", -- 7 
					"0000000" when "00001000", -- 8
					"0001100" when "00001001", -- 9
					--Letters/repeat-----------
					"0000001" when "00001010", -- 0
					"1001111" when "00001011", -- 1
					"0010010" when "00001100", -- 2
					"0000110" when "00001101", -- 3
				   "1001100" when "00001110", -- 4
			      "0100100" when "00001111", -- 5
					"0100000" when "00010000", -- 6
					"0001111" when "00010001", -- 7
					"0000000" when "00010010", -- 8
					"0001100" when "00010011", -- 9
					
					"0000001" when "00010100", -- 0
					"1001111" when "00010101", -- 1
					"0010010" when "00010110", -- 2
					"0000110" when "00010111", -- 3
					"1001100" when "00011000", -- 4
					"0100100" when "00011001", -- 5
					"0100000" when "00011010", -- 6
					"0001111" when "00011011", -- 7
					"0000000" when "00011100", -- 8
					"0001100" when "00011101", -- 9
					
					"0000001" when "00011110", -- 0
					"1001111" when "00011111", -- 1
					"0010010" when "00100000", -- 2
					"0000110" when "00100001", -- 3
					"1001100" when "00100010", -- 4
					"0100100" when "00100011", -- 5
					"0100000" when "00100100", -- 6
					"0001111" when "00100101", -- 7
					"0000000" when "00100110", -- 8
					"0001100" when "00100111", -- 9
					
					"0000001" when "00101000", -- 0
					"1001111" when "00101001", -- 1
					"0010010" when "00101010", -- 2
					"0000110" when "00101011", -- 3
					"1001100" when "00101100", -- 4
					"0100100" when "00101101", -- 5
					"0100000" when "00101110", -- 6
					"0001111" when "00101111", -- 7
					"0000000" when "00110000", -- 8
					"0001100" when "00110001", -- 9
					
					"0000001" when "00110010", -- 0
					
					"1111111" when others;
					
					
					-------------------------------------------------------------------
  with (SW) select 
  HEX1 <= "0000001" when "00000000", -- 0
               "0000001" when "00000001", -- 0
					"0000001" when "00000010", -- 0
					"0000001" when "00000011", -- 0
					"0000001" when "00000100", -- 0
					"0000001" when "00000101", -- 0
					"0000001" when "00000110", -- 0 
					"0000001" when "00000111", -- 0 
					"0000001" when "00001000", -- 0
					"0000001" when "00001001", -- 0
					
					"1001111" when "00001010", -- 1
					"1001111" when "00001011", -- 1
					"1001111" when "00001100", -- 1
					"1001111" when "00001101", -- 1
				   "1001111" when "00001110", -- 1
			      "1001111" when "00001111", -- 1
					"1001111" when "00010000", -- 1
					"1001111" when "00010001", -- 1
					"1001111" when "00010010", -- 1
					"1001111" when "00010011", -- 1
					
					"0010010" when "00010100", -- 2
					"0010010" when "00010101", -- 2
					"0010010" when "00010110", -- 2
					"0010010" when "00010111", -- 2
					"0010010" when "00011000", -- 2
					"0010010" when "00011001", -- 2
					"0010010" when "00011010", -- 2
					"0010010" when "00011011", -- 2
					"0010010" when "00011100", -- 2
					"0010010" when "00011101", -- 2
					
					"0000110" when "00011110", -- 3
					"0000110" when "00011111", -- 3
					"0000110" when "00100000", -- 3
					"0000110" when "00100001", -- 3
					"0000110" when "00100010", -- 3
					"0000110" when "00100011", -- 3
					"0000110" when "00100100", -- 3
					"0000110" when "00100101", -- 3
					"0000110" when "00100110", -- 3
					"0000110" when "00100111", -- 3
					
					"1001100" when "00101000", -- 4
					"1001100" when "00101001", -- 4
					"1001100" when "00101010", -- 4
					"1001100" when "00101011", -- 4
					"1001100" when "00101100", -- 4
					"1001100" when "00101101", -- 4
					"1001100" when "00101110", -- 4
					"1001100" when "00101111", -- 4
					"1001100" when "00110000", -- 4
					"1001100" when "00110001", -- 4
					
					"0100100" when "00110010", -- 5
					
					"1111111" when others;
					

end decoder_arch; 